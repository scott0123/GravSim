//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Changed the purpose of this file. Now must return is_ball based on --
//        inputted position of ball.												 --
//-------------------------------------------------------------------------


module  ball ( input         Clk,                // 50 MHz clock
                             Reset,              // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
//               input [7:0]   keycode,            // Keycode from the keyboard
               input [9:0]   DrawX, DrawY,       // Current pixel coordinates
					
					input [31:0]  radius, posX, posY, posZ,
					
               output logic  is_ball             // Whether current pixel belongs to ball or background
              );
    
    parameter [9:0] Ball_X_Center = 10'd320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center = 10'd240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min = 10'd0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max = 10'd639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min = 10'd0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max = 10'd479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step = 10'd1;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step = 10'd1;      // Step size on the Y axis
    parameter [9:0] Ball_Size = 10'd4;        // Ball size

//    parameter [7:0] KEYCODE_UP = 8'd26;                  // Keycode for the key UP (in this case: W)
//    parameter [7:0] KEYCODE_DOWN = 8'd22;                  // Keycode for the key DOWN (in this case: S)
//    parameter [7:0] KEYCODE_LEFT = 8'd4;                  // Keycode for the key LEFT (in this case: A)
//    parameter [7:0] KEYCODE_RIGHT = 8'd7;                  // Keycode for the key RIGHT (in this case: D)
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
    logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
    
    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    //////// Do not modify the always_ff blocks. ////////
    
    // Compute whether the pixel corresponds to ball or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
    int DistX, DistY, Size;
    assign DistX = DrawX - posX;
    assign DistY = DrawY - posY;
	 
	 // absolute value of Dists
	 int absDistX, absDistY;
	 
	 logic [31:0] adjRadius;

	 // perform absolute value operations and calculate Z size adjust limit
	 always_comb begin
//		if ( DistX < 0 ) begin
//			absDistX = -DistX;
//		end
//		else begin
//			absDistX = DistX;
//		end
//		
//		if ( DistY < 0 ) begin
//			absDistY = -DistY;
//		end
//		else begin
//			absDistY = DistY;
//		end
		
		// radius adjust
		if ( posZ < 1 ) begin
			adjRadius = 1;
		end
		else if ( posZ > 80 ) begin
			adjRadius = 80;
		end
		else begin
			adjRadius = posZ;
		end
		
	 end
	 
	 // currently depends ONLY on Z
    assign Size = adjRadius;
	 
    always_comb begin
        if ( ( DistX*DistX + DistY*DistY) <= (Size*Size) )
//			if ( ( absDistX + absDistY) <= (Size) )
            is_ball = 1'b1;
        else
            is_ball = 1'b0;
        /* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while 
           the single line is quite powerful descriptively, it causes the synthesis tool to use up three
           of the 12 available multipliers on the chip! */
    end
    
endmodule
