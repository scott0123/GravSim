//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Changed the purpose of this file. Now must return is_ball based on --
//        inputted position of ball.												 --
//-------------------------------------------------------------------------


module  ball ( input         Clk,                // 50 MHz clock
                             Reset,              // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
//               input [7:0]   keycode,            // Keycode from the keyboard
               input [9:0]   DrawX, DrawY,       // Current pixel coordinates
					
					input [31:0]  radius, posX, posY, posZ, // floats
					
               output logic  is_ball             // Whether current pixel belongs to ball or background
              );
    
	 // consts needed to scale radius, posX, posY, posZ
	 const int FLOAT2 = 32'h40000000;
	 const int FLOAT10 = 32'h41200000;
	 const int FLOAT100 = 32'h42c80000;
	 
	 
    parameter [9:0] Ball_X_Center = 10'd320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center = 10'd240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min = 10'd0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max = 10'd639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min = 10'd0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max = 10'd479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step = 10'd1;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step = 10'd1;      // Step size on the Y axis
    parameter [9:0] Ball_Size = 10'd4;        // Ball size

//    parameter [7:0] KEYCODE_UP = 8'd26;                  // Keycode for the key UP (in this case: W)
//    parameter [7:0] KEYCODE_DOWN = 8'd22;                  // Keycode for the key DOWN (in this case: S)
//    parameter [7:0] KEYCODE_LEFT = 8'd4;                  // Keycode for the key LEFT (in this case: A)
//    parameter [7:0] KEYCODE_RIGHT = 8'd7;                  // Keycode for the key RIGHT (in this case: D)
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
    logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
    
	 // integer (pixel) versions of radius, posX, posY, posZ
	 logic [31:0] intRad, intPosX, intPosY, intPosZ;
	 
	 always_comb begin
	 
		
	 
	 end
	 
	 
	 
    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    //////// Do not modify the always_ff blocks. ////////
    
    // Compute whether the pixel corresponds to ball or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
    int DistX, DistY, Size;
    assign DistX = DrawX - (intPosX + 32'd320);
    assign DistY = DrawY - (intPosY + 32'd240);
	 
	 // absolute value of Dists
	 int absDistX, absDistY;
	 
	 logic [31:0] adjRadius;

	 // perform absolute value operations and calculate Z size adjust limit
	 always_comb begin
		
		// radius adjust
		if ( (intPosZ + 32'd20) < 1 ) begin
			adjRadius = 1;
		end
		else if ( (intPosZ + 32'd20) > 80 ) begin
			adjRadius = 80;
		end
		else begin
			adjRadius = (intPosZ + 32'd20);
		end
		
	 end
	 
	 // currently depends ONLY on Z
    assign Size = adjRadius;
	 
    always_comb begin
        if ( ( DistX*DistX + DistY*DistY) <= (Size*Size) )
//			if ( ( absDistX + absDistY) <= (Size) )
            is_ball = 1'b1;
        else
            is_ball = 1'b0;
        /* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while 
           the single line is quite powerful descriptively, it causes the synthesis tool to use up three
           of the 12 available multipliers on the chip! */
    end



// -----------------------------------------------------------------

//	   Modules are instantiated here so they have access to regfile

// -----------------------------------------------------------------


logic [31:0] FPmultRad_out;
logic [31:0] FPmultX_out;
logic [31:0] FPmultY_out;
logic [31:0] FPmultZ_out;
logic [31:0] FPaddX_out;
logic [31:0] FPaddY_out;
logic [31:0] FPaddZ_out;

FPmult FPmultRad (
	// inputs
	.iA(radius),
	.iB(FLOAT10),
	// outputs
	.oProd(FPmultRad_out)
);

FPmult FPmultX (
	// inputs
	.iA(posX),
	.iB(FLOAT100),
	// outputs
	.oProd(FPmultX_out)
);

FPmult FPmultY (
	// inputs
	.iA(posY),
	.iB(FLOAT100),
	// outputs
	.oProd(FPmultY_out)
);

FPmult FPmultZ (
	// inputs
	.iA(posZ),
	.iB(FLOAT2),
	// outputs
	.oProd(FPmultZ_out)
);

fp2int fp2intRad (
	// inputs
	.fp_in(FPmultRad_out),
	//outputs
	.int_out(intRad)
);

fp2int fp2intX (
	// inputs
	.fp_in(FPmultX_out),
	//outputs
	.int_out(intPosX)
);

fp2int fp2intY (
	// inputs
	.fp_in(FPmultY_out),
	//outputs
	.int_out(intPosY)
);

fp2int fp2intZ (
	// inputs
	.fp_in(FPmultZ_out),
	//outputs
	.int_out(intPosZ)
);

endmodule
